class fa_sqr extends uvm_sequencer #(fa_tran);
  `uvm_component_utils(fa_sqr)

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction
endclass
