class spi_drv extends uvm_driver #(spi_tran);
  `uvm_component_utils(spi_drv)

  virtual spi_if vif;
  uvm_analysis_port #(spi_tran) drv_ap;

  function new(string name, uvm_component parent);
    super.new(name, parent);
    drv_ap = new("drv_ap", this);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if(!uvm_config_db#(virtual spi_if)::get(this, "", "vif", vif)) begin
      `uvm_error("DRIVER", "Virtual interface (spi_if) not found in config db")
    end
  endfunction

  task run_phase(uvm_phase phase);
    spi_tran tr;
    forever begin
      seq_item_port.get_next_item(tr);
//
      @(vif.drv_cb);
	`uvm_info(get_type_name(), "Good news for seeing this", UVM_LOW)
//      uvm_config_db#(int)::set(null, "*", "tran_count", tr.seq_count);
//      uvm_config_db#(int)::set(null, "*", "tran_index", tr.seq_index);
//      uvm_config_db#(string)::set(null, "*", "tran_type", tr.seq_type);
//
//      `uvm_info("DRIVER", $sformatf("Drive %0d/%0d %s tran to DUT: a=%0b, b=%0b, cin=%0b",
//                                    tr.seq_index, tr.seq_count, tr.seq_type, tr.a, tr.b, tr.cin),
//                                    UVM_MEDIUM)
//
//      vif.drv_cb.a_tb   <= tr.a;      // Drive 'a' from transaction (tr) to DUT
//      vif.drv_cb.b_tb   <= tr.b;      // Drive 'b' from transaction (tr) to DUT
//      vif.drv_cb.cin_tb <= tr.cin;  // Drive 'cin' from transaction (tr) to DUT
//
      seq_item_port.item_done();
    end
  endtask
endclass

