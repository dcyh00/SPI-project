`include "spi_test.sv"
`include "spi_protocol_test.sv"
`include "spi_start_test.sv"
