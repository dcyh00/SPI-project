`include "spi_seq.sv"
`include "protocol_seq.sv"
`include "random_seq.sv"
