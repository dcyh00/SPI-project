`include "spi_seq.sv"
`include "protocol_seq.sv"
